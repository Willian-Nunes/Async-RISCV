/*/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////// BYPASS UNIT ////////////////////////////////////////////////////////////////
 //////////////////////////////////////// Developed By: Willian Analdo Nunes ///////////////////////////////////////////////////
 //////////////////////////////////////////// PUCRS, Porto Alegre, 2020      ///////////////////////////////////////////////////
 /////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////*/

`include "pkg.sv"
import my_pkg::*;

module bypassUnit #(parameter  DEPTH = 3)           // LUI, NOP E INVALID
    (input logic clk,
    input logic [31:0]  opA,
    output logic [31:0] result_out);

    logic [31:0] result[DEPTH];

    assign result_out = result[DEPTH-1];

    always @(posedge clk) begin
        result[0] <= opA;
        
        for(int i = 1; i < DEPTH; i++)
            result[i] <= result[i-1];
    end
endmodule

